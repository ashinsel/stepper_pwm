library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package config is
end package;

package body config is
end config;


